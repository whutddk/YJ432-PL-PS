//////////////////////////////////////////////////////////////////////////////////
// Company:   
// Engineer: Ruige_Lee
// Create Date: 2019-05-24 14:15:27
// Last Modified by:   Ruige_Lee
// Last Modified time: 2019-05-24 14:22:05
// Email: 295054118@whut.edu.cn
// page: https://whutddk.github.io/
// Design Name:   
// Module Name: PartialReconfigurationTop
// Project Name:   
// Target Devices:   
// Tool Versions:   
// Description:   
// 
// Dependencies:   
// 
// Revision:  
// Revision:    -   
// Additional Comments:  
// 
//
//////////////////////////////////////////////////////////////////////////////////


module PartialReconfigurationTop (
	input CLK,
	input RST_n,
	



);





endmodule


