//////////////////////////////////////////////////////////////////////////////////
// Company: WUT  
// Engineer: WUT RUIGE LEE
// Create Date: 2018/06/21 10:07:43
// Last Modified by:   WUT_Ruige_Lee
// Last Modified time: 2019-01-12 16:39:00
// Email: 295054118@whut.edu.cn
// Design Name:   
// Module Name: ip_SRAM
// Project Name:   
// Target Devices:   
// Tool Versions:   
// Description:   
// 
// Dependencies:   
// 
// Revision:  
// Revision 0.01 - File Created
// Additional Comments:  
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps


module perip_SRAM(    
);
	
	
endmodule
