//////////////////////////////////////////////////////////////////////////////////
// Company:  WUT
// Engineer: WUT RUIGE LEE
// Create Date: 2018/06/21 17:44:39
// Last Modified by:   WUT_Ruige_Lee
// Last Modified time: 2019-01-12 16:16:26
// Email: 295054118@whut.edu.cn
// Design Name:   
// Module Name: FB_SWKEY
// Project Name:   
// Target Devices:   
// Tool Versions:   
// Description:   
// 
// Dependencies:   
// 
// Revision:  
// Revision 0.01 - File Created
// Additional Comments:  
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps


module FB_SWKEY(
	
    );
endmodule